library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity onetofourdemuxwithenable is
    Port ( );
end onetofourdemuxwithenable;

architecture Behavioral of onetofourdemuxwithenable is

begin


end Behavioral;
