library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity fourtoonebusmux is
    Port ( );
end fourtoonebusmux;

architecture Behavioral of fourtoonebusmux is

begin


end Behavioral;
